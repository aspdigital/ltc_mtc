-------------------------------------------------------------------------------
-- Title      : Choose what to display on the 7-segment LEDs
-- Project    : 
-------------------------------------------------------------------------------
-- File       : display_mux.vhdl
-- Author     : Andy Peters  <devel@latke.net>
-- Company    : ASP Digital
-- Created    : 2025-05-12
-- Last update: 2025-05-12
-- Platform   : 
-- Standard   : VHDL'08, Math Packages
-------------------------------------------------------------------------------
-- Description: There are three things that can drive the LED timecode display.
-- They are:
-- 1. The time code generator, which also feeds both the LTC and MTC outputs,
-- 2. The MTC receiver,
-- 3. The LTC receiver.
--
-- Two switches determine what is displayed:
-- a. Internal/External,
-- b. MTC/LTC if in external mode.
--
-- The three sources have the time code and the frame rate. Based on the source selects and the chosen frame
-- rate, we choose the timer clock. The selected time code is synchronized to that clock and that's what
-- drives the display logic.
-------------------------------------------------------------------------------
-- Copyright (c) 2025 ASP Digital
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2025-05-12  -        andy    Created
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity display_mux is
    generic (
        CLKPER_30FPS : time;
        CLKPER_25FPS : time;
        CLKPER_24FPS : time);
    port (
        -- main clock, for selection
        clk_main        : in  std_logic;
        rst_main        : in  std_logic;
        -- so we know we have timer clocks.
        mmcm_locked     : in  std_logic;
        -- all of the timer clocks.
        clk_bundle      : in  clk_bundle_t;
        -- display select.
        tc_display_src  : in std_logic;  -- 0 = internal, 1 = external
        tc_ext_src      : in std_logic;  -- 0 = mtc, 1 = ltcXS
        -- the frame rate and time generated by the local timer
        gen_frame_time  : in  frame_time_t;
        gen_frame_rate  : in  frame_rate_t;
        -- decoded frame rate and time received from the MIDI port.
        mtcd_frame_time : in  frame_time_t;
        mtcd_frame_rate : in  frame_rate_t;
        -- decode frame rate and time received from the LTC in port.
        ltcd_frame_time : in  frame_time_t;
        ltcd_frame_rate : in  frame_rate_t;
        -- all of the LED segments to display the current selected time code
        display         : out display_t);
end entity display_mux;

architecture mux of display_mux is

    -- frame rate based on the selects.

begin  -- architecture mux

    -- timer clock frequency is determined by the selected frame rate.
    display_clk_mux : entity work.clk_mux(mux)
        port map (
            clk_main    => clk_main,
            rst_main    => rst_main,
            mmcm_locked => mmcm_locked,
            frame_rate  => frame_rate,
            clk_bundle  => clk_bundle,
            clk_out     => clk_out,
            rst_out     => rst_out);
    
    tcd : entity work.timecode_display(digit_driver)
        generic map (
            CLKPER_30FPS => CLKPER_30FPS,
            CLKPER_25FPS => CLKPER_25FPS,
            CLKPER_24FPS => CLKPER_24FPS)
        port map (
            clk_timer  => clk_timer,
            rst_timer  => rst_timer,
            frame_time => frame_time,
            frame_rate => frame_rate_s,
            display    => display);

end architecture mux;
