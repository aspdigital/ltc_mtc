-------------------------------------------------------------------------------
-- Title      : Linear Time Code Decoder
-- Project    : 
-------------------------------------------------------------------------------
-- File       : ltc_decode.vhdl
-- Author     : Andy Peters  <devel@latke.net>
-- Company    : ASP Digital
-- Created    : 2025-04-20
-- Last update: 2025-05-14
-- Platform   : 
-- Standard   : VHDL'08, Math Packages
-------------------------------------------------------------------------------
-- Description: Decode the incoming time code.
-------------------------------------------------------------------------------
-- Copyright (c) 2025 ASP Digital
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2025-04-20  -        andy	Created
-------------------------------------------------------------------------------
entity ltc_decode is
  
end entity ltc_decode;

architecture decoder of ltc_decode is

begin  -- architecture decoder

  

end architecture decoder;



